library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

Entity MemoriaROM16bits is 
	Port
	(
		adress: in unsigned(4 downto 0);
		enable: in std_logic;
		saida: out unsigned(15 downto 0)
	);
End MemoriaROM16bits;

Architecture behavior of MemoriaROM16bits is

	Type pattern is array (Natural Range <>) of unsigned(15 downto 0);
	
	constant data : pattern (0 to 31):=
	
	(
"0000000000000000","0000000000000001","0000000000000010","0000000000000011", "0000000000000100","0000000000000101","0000000000000110","0000000000000111",
					 
"0000000000001000","0000000000001001","0000000000001010","0000000000001011", "0000000000001100","0000000000001101","0000000000001110","0000000000001111",
					 
"0000000000010000","0000000000010001","0000000000010010","0000000000010011", "0000000000010100","0000000000010101","0000000000010110","0000000000010111",
					 
"0000000000011000","0000000000011001","0000000000011010","0000000000011011", "0000000000011100","0000000000011101","0000000000011110","0000000000011111"  );

	BEGIN
		
		saida <= data(to_integer(adress)) when enable='0' else (Others=>'Z');
		
	End behavior;