LIBRARY ieee; USE ieee.std_logic_1164.all; USE ieee.numeric_std.all; USE ieee.std_logic_unsigned.all;

ENTITY MemoriaRAM16bits IS
 PORT(
		ADDRESS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		DATA : INOUT STD_LOGIC_VECTOR (3 DOWNTO 0); 
		WR : IN STD_LOGIC; 
		RD : IN STD_LOGIC 
 );

END ENTITY;

ARCHITECTURE COMPORTAMENTO OF MemoriaRAM16bits IS

	TYPE RAM IS ARRAY (INTEGER RANGE <>) OF STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL DATA_OUT : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL MEM : RAM (0 TO 15);

BEGIN
 --TRI-STATE BUFFER CONTROL (N ENTENDI ESSA PARTE)
 DATA <= DATA_OUT WHEN (RD = '1') ELSE (OTHERS => 'Z');
 
 MEM_WRITE: PROCESS(ADDRESS, DATA, WR)
	BEGIN
		IF (WR = '1') THEN
		
			MEM(TO_INTEGER(UNSIGNED(ADDRESS))) <= DATA;
			
		END IF;
	END PROCESS;

 MEM_READ: PROCESS(ADDRESS, RD)
	BEGIN
		IF(RD = '1') THEN
		
			DATA_OUT <= MEM(TO_INTEGER(UNSIGNED(ADDRESS)));
			
		END IF;
	END PROCESS;
	
END ARCHITECTURE;  
